
* .GLOBAL VDD! GND

.subckt CIM_arr in0 in1 in2 in3 in4 in5 in6 in7 in8 in9
+ in10 in11 in12 in13 in14 in15 in16 in17 in18 in19
+ in20 in21 in22 in23 in24 in25 in26 in27 in28 in29
+ in30 in31
+ Prod0_0[3] Prod0_0[2] Prod0_0[1] Prod0_0[0]
+ Prod0_1[3] Prod0_1[2] Prod0_1[1] Prod0_1[0]
+ Prod0_2[3] Prod0_2[2] Prod0_2[1] Prod0_2[0]
+ Prod0_3[3] Prod0_3[2] Prod0_3[1] Prod0_3[0]
+ Prod0_4[3] Prod0_4[2] Prod0_4[1] Prod0_4[0]
+ Prod0_5[3] Prod0_5[2] Prod0_5[1] Prod0_5[0]
+ Prod0_6[3] Prod0_6[2] Prod0_6[1] Prod0_6[0]
+ Prod0_7[3] Prod0_7[2] Prod0_7[1] Prod0_7[0]
+ Prod0_8[3] Prod0_8[2] Prod0_8[1] Prod0_8[0]
+ Prod0_9[3] Prod0_9[2] Prod0_9[1] Prod0_9[0]
+ Prod0_10[3] Prod0_10[2] Prod0_10[1] Prod0_10[0]
+ Prod0_11[3] Prod0_11[2] Prod0_11[1] Prod0_11[0]
+ Prod0_12[3] Prod0_12[2] Prod0_12[1] Prod0_12[0]
+ Prod0_13[3] Prod0_13[2] Prod0_13[1] Prod0_13[0]
+ Prod0_14[3] Prod0_14[2] Prod0_14[1] Prod0_14[0]
+ Prod0_15[3] Prod0_15[2] Prod0_15[1] Prod0_15[0]
+ Prod0_16[3] Prod0_16[2] Prod0_16[1] Prod0_16[0]
+ Prod0_17[3] Prod0_17[2] Prod0_17[1] Prod0_17[0]
+ Prod0_18[3] Prod0_18[2] Prod0_18[1] Prod0_18[0]
+ Prod0_19[3] Prod0_19[2] Prod0_19[1] Prod0_19[0]
+ Prod0_20[3] Prod0_20[2] Prod0_20[1] Prod0_20[0]
+ Prod0_21[3] Prod0_21[2] Prod0_21[1] Prod0_21[0]
+ Prod0_22[3] Prod0_22[2] Prod0_22[1] Prod0_22[0]
+ Prod0_23[3] Prod0_23[2] Prod0_23[1] Prod0_23[0]
+ Prod0_24[3] Prod0_24[2] Prod0_24[1] Prod0_24[0]
+ Prod0_25[3] Prod0_25[2] Prod0_25[1] Prod0_25[0]
+ Prod0_26[3] Prod0_26[2] Prod0_26[1] Prod0_26[0]
+ Prod0_27[3] Prod0_27[2] Prod0_27[1] Prod0_27[0]
+ Prod0_28[3] Prod0_28[2] Prod0_28[1] Prod0_28[0]
+ Prod0_29[3] Prod0_29[2] Prod0_29[1] Prod0_29[0]
+ Prod0_30[3] Prod0_30[2] Prod0_30[1] Prod0_30[0]
+ Prod0_31[3] Prod0_31[2] Prod0_31[1] Prod0_31[0]
+ Prod1_0[3] Prod1_0[2] Prod1_0[1] Prod1_0[0]
+ Prod1_1[3] Prod1_1[2] Prod1_1[1] Prod1_1[0]
+ Prod1_2[3] Prod1_2[2] Prod1_2[1] Prod1_2[0]
+ Prod1_3[3] Prod1_3[2] Prod1_3[1] Prod1_3[0]
+ Prod1_4[3] Prod1_4[2] Prod1_4[1] Prod1_4[0]
+ Prod1_5[3] Prod1_5[2] Prod1_5[1] Prod1_5[0]
+ Prod1_6[3] Prod1_6[2] Prod1_6[1] Prod1_6[0]
+ Prod1_7[3] Prod1_7[2] Prod1_7[1] Prod1_7[0]
+ Prod1_8[3] Prod1_8[2] Prod1_8[1] Prod1_8[0]
+ Prod1_9[3] Prod1_9[2] Prod1_9[1] Prod1_9[0]
+ Prod1_10[3] Prod1_10[2] Prod1_10[1] Prod1_10[0]
+ Prod1_11[3] Prod1_11[2] Prod1_11[1] Prod1_11[0]
+ Prod1_12[3] Prod1_12[2] Prod1_12[1] Prod1_12[0]
+ Prod1_13[3] Prod1_13[2] Prod1_13[1] Prod1_13[0]
+ Prod1_14[3] Prod1_14[2] Prod1_14[1] Prod1_14[0]
+ Prod1_15[3] Prod1_15[2] Prod1_15[1] Prod1_15[0]
+ Prod1_16[3] Prod1_16[2] Prod1_16[1] Prod1_16[0]
+ Prod1_17[3] Prod1_17[2] Prod1_17[1] Prod1_17[0]
+ Prod1_18[3] Prod1_18[2] Prod1_18[1] Prod1_18[0]
+ Prod1_19[3] Prod1_19[2] Prod1_19[1] Prod1_19[0]
+ Prod1_20[3] Prod1_20[2] Prod1_20[1] Prod1_20[0]
+ Prod1_21[3] Prod1_21[2] Prod1_21[1] Prod1_21[0]
+ Prod1_22[3] Prod1_22[2] Prod1_22[1] Prod1_22[0]
+ Prod1_23[3] Prod1_23[2] Prod1_23[1] Prod1_23[0]
+ Prod1_24[3] Prod1_24[2] Prod1_24[1] Prod1_24[0]
+ Prod1_25[3] Prod1_25[2] Prod1_25[1] Prod1_25[0]
+ Prod1_26[3] Prod1_26[2] Prod1_26[1] Prod1_26[0]
+ Prod1_27[3] Prod1_27[2] Prod1_27[1] Prod1_27[0]
+ Prod1_28[3] Prod1_28[2] Prod1_28[1] Prod1_28[0]
+ Prod1_29[3] Prod1_29[2] Prod1_29[1] Prod1_29[0]
+ Prod1_30[3] Prod1_30[2] Prod1_30[1] Prod1_30[0]
+ Prod1_31[3] Prod1_31[2] Prod1_31[1] Prod1_31[0]
+ Prod2_0[3] Prod2_0[2] Prod2_0[1] Prod2_0[0]
+ Prod2_1[3] Prod2_1[2] Prod2_1[1] Prod2_1[0]
+ Prod2_2[3] Prod2_2[2] Prod2_2[1] Prod2_2[0]
+ Prod2_3[3] Prod2_3[2] Prod2_3[1] Prod2_3[0]
+ Prod2_4[3] Prod2_4[2] Prod2_4[1] Prod2_4[0]
+ Prod2_5[3] Prod2_5[2] Prod2_5[1] Prod2_5[0]
+ Prod2_6[3] Prod2_6[2] Prod2_6[1] Prod2_6[0]
+ Prod2_7[3] Prod2_7[2] Prod2_7[1] Prod2_7[0]
+ Prod2_8[3] Prod2_8[2] Prod2_8[1] Prod2_8[0]
+ Prod2_9[3] Prod2_9[2] Prod2_9[1] Prod2_9[0]
+ Prod2_10[3] Prod2_10[2] Prod2_10[1] Prod2_10[0]
+ Prod2_11[3] Prod2_11[2] Prod2_11[1] Prod2_11[0]
+ Prod2_12[3] Prod2_12[2] Prod2_12[1] Prod2_12[0]
+ Prod2_13[3] Prod2_13[2] Prod2_13[1] Prod2_13[0]
+ Prod2_14[3] Prod2_14[2] Prod2_14[1] Prod2_14[0]
+ Prod2_15[3] Prod2_15[2] Prod2_15[1] Prod2_15[0]
+ Prod2_16[3] Prod2_16[2] Prod2_16[1] Prod2_16[0]
+ Prod2_17[3] Prod2_17[2] Prod2_17[1] Prod2_17[0]
+ Prod2_18[3] Prod2_18[2] Prod2_18[1] Prod2_18[0]
+ Prod2_19[3] Prod2_19[2] Prod2_19[1] Prod2_19[0]
+ Prod2_20[3] Prod2_20[2] Prod2_20[1] Prod2_20[0]
+ Prod2_21[3] Prod2_21[2] Prod2_21[1] Prod2_21[0]
+ Prod2_22[3] Prod2_22[2] Prod2_22[1] Prod2_22[0]
+ Prod2_23[3] Prod2_23[2] Prod2_23[1] Prod2_23[0]
+ Prod2_24[3] Prod2_24[2] Prod2_24[1] Prod2_24[0]
+ Prod2_25[3] Prod2_25[2] Prod2_25[1] Prod2_25[0]
+ Prod2_26[3] Prod2_26[2] Prod2_26[1] Prod2_26[0]
+ Prod2_27[3] Prod2_27[2] Prod2_27[1] Prod2_27[0]
+ Prod2_28[3] Prod2_28[2] Prod2_28[1] Prod2_28[0]
+ Prod2_29[3] Prod2_29[2] Prod2_29[1] Prod2_29[0]
+ Prod2_30[3] Prod2_30[2] Prod2_30[1] Prod2_30[0]
+ Prod2_31[3] Prod2_31[2] Prod2_31[1] Prod2_31[0]
+ Prod3_0[3] Prod3_0[2] Prod3_0[1] Prod3_0[0]
+ Prod3_1[3] Prod3_1[2] Prod3_1[1] Prod3_1[0]
+ Prod3_2[3] Prod3_2[2] Prod3_2[1] Prod3_2[0]
+ Prod3_3[3] Prod3_3[2] Prod3_3[1] Prod3_3[0]
+ Prod3_4[3] Prod3_4[2] Prod3_4[1] Prod3_4[0]
+ Prod3_5[3] Prod3_5[2] Prod3_5[1] Prod3_5[0]
+ Prod3_6[3] Prod3_6[2] Prod3_6[1] Prod3_6[0]
+ Prod3_7[3] Prod3_7[2] Prod3_7[1] Prod3_7[0]
+ Prod3_8[3] Prod3_8[2] Prod3_8[1] Prod3_8[0]
+ Prod3_9[3] Prod3_9[2] Prod3_9[1] Prod3_9[0]
+ Prod3_10[3] Prod3_10[2] Prod3_10[1] Prod3_10[0]
+ Prod3_11[3] Prod3_11[2] Prod3_11[1] Prod3_11[0]
+ Prod3_12[3] Prod3_12[2] Prod3_12[1] Prod3_12[0]
+ Prod3_13[3] Prod3_13[2] Prod3_13[1] Prod3_13[0]
+ Prod3_14[3] Prod3_14[2] Prod3_14[1] Prod3_14[0]
+ Prod3_15[3] Prod3_15[2] Prod3_15[1] Prod3_15[0]
+ Prod3_16[3] Prod3_16[2] Prod3_16[1] Prod3_16[0]
+ Prod3_17[3] Prod3_17[2] Prod3_17[1] Prod3_17[0]
+ Prod3_18[3] Prod3_18[2] Prod3_18[1] Prod3_18[0]
+ Prod3_19[3] Prod3_19[2] Prod3_19[1] Prod3_19[0]
+ Prod3_20[3] Prod3_20[2] Prod3_20[1] Prod3_20[0]
+ Prod3_21[3] Prod3_21[2] Prod3_21[1] Prod3_21[0]
+ Prod3_22[3] Prod3_22[2] Prod3_22[1] Prod3_22[0]
+ Prod3_23[3] Prod3_23[2] Prod3_23[1] Prod3_23[0]
+ Prod3_24[3] Prod3_24[2] Prod3_24[1] Prod3_24[0]
+ Prod3_25[3] Prod3_25[2] Prod3_25[1] Prod3_25[0]
+ Prod3_26[3] Prod3_26[2] Prod3_26[1] Prod3_26[0]
+ Prod3_27[3] Prod3_27[2] Prod3_27[1] Prod3_27[0]
+ Prod3_28[3] Prod3_28[2] Prod3_28[1] Prod3_28[0]
+ Prod3_29[3] Prod3_29[2] Prod3_29[1] Prod3_29[0]
+ Prod3_30[3] Prod3_30[2] Prod3_30[1] Prod3_30[0]
+ Prod3_31[3] Prod3_31[2] Prod3_31[1] Prod3_31[0]

X_inv0 in0 VDD! GND in0_b INVx13_ASAP7_75t_R 
X_inv1 in1 VDD! GND in1_b INVx13_ASAP7_75t_R 
X_inv2 in2 VDD! GND in2_b INVx13_ASAP7_75t_R 
X_inv3 in3 VDD! GND in3_b INVx13_ASAP7_75t_R 
X_inv4 in4 VDD! GND in4_b INVx13_ASAP7_75t_R 
X_inv5 in5 VDD! GND in5_b INVx13_ASAP7_75t_R 
X_inv6 in6 VDD! GND in6_b INVx13_ASAP7_75t_R 
X_inv7 in7 VDD! GND in7_b INVx13_ASAP7_75t_R 
X_inv8 in8 VDD! GND in8_b INVx13_ASAP7_75t_R 
X_inv9 in9 VDD! GND in9_b INVx13_ASAP7_75t_R 

X_inv10 in10 VDD! GND in10_b INVx13_ASAP7_75t_R 
X_inv11 in11 VDD! GND in11_b INVx13_ASAP7_75t_R 
X_inv12 in12 VDD! GND in12_b INVx13_ASAP7_75t_R 
X_inv13 in13 VDD! GND in13_b INVx13_ASAP7_75t_R 
X_inv14 in14 VDD! GND in14_b INVx13_ASAP7_75t_R 
X_inv15 in15 VDD! GND in15_b INVx13_ASAP7_75t_R 
X_inv16 in16 VDD! GND in16_b INVx13_ASAP7_75t_R 
X_inv17 in17 VDD! GND in17_b INVx13_ASAP7_75t_R 
X_inv18 in18 VDD! GND in18_b INVx13_ASAP7_75t_R 
X_inv19 in19 VDD! GND in19_b INVx13_ASAP7_75t_R 
                      
X_inv20 in20 VDD! GND in20_b INVx13_ASAP7_75t_R 
X_inv21 in21 VDD! GND in21_b INVx13_ASAP7_75t_R 
X_inv22 in22 VDD! GND in22_b INVx13_ASAP7_75t_R 
X_inv23 in23 VDD! GND in23_b INVx13_ASAP7_75t_R 
X_inv24 in24 VDD! GND in24_b INVx13_ASAP7_75t_R 
X_inv25 in25 VDD! GND in25_b INVx13_ASAP7_75t_R 
X_inv26 in26 VDD! GND in26_b INVx13_ASAP7_75t_R 
X_inv27 in27 VDD! GND in27_b INVx13_ASAP7_75t_R 
X_inv28 in28 VDD! GND in28_b INVx13_ASAP7_75t_R 
X_inv29 in29 VDD! GND in29_b INVx13_ASAP7_75t_R 
                      
X_inv30 in30 VDD! GND in30_b INVx13_ASAP7_75t_R 
X_inv31 in31 VDD! GND in31_b INVx13_ASAP7_75t_R 

X_Wcol0 in0_b in1_b in2_b in3_b in4_b in5_b in6_b in7_b in8_b in9_b
+ in10_b in11_b in12_b in13_b in14_b in15_b in16_b in17_b in18_b in19_b
+ in20_b in21_b in22_b in23_b in24_b in25_b in26_b in27_b in28_b in29_b
+ in30_b in31_b
+ Prod0_0[3] Prod0_0[2] Prod0_0[1] Prod0_0[0]
+ Prod0_1[3] Prod0_1[2] Prod0_1[1] Prod0_1[0]
+ Prod0_2[3] Prod0_2[2] Prod0_2[1] Prod0_2[0]
+ Prod0_3[3] Prod0_3[2] Prod0_3[1] Prod0_3[0]
+ Prod0_4[3] Prod0_4[2] Prod0_4[1] Prod0_4[0]
+ Prod0_5[3] Prod0_5[2] Prod0_5[1] Prod0_5[0]
+ Prod0_6[3] Prod0_6[2] Prod0_6[1] Prod0_6[0]
+ Prod0_7[3] Prod0_7[2] Prod0_7[1] Prod0_7[0]
+ Prod0_8[3] Prod0_8[2] Prod0_8[1] Prod0_8[0]
+ Prod0_9[3] Prod0_9[2] Prod0_9[1] Prod0_9[0]
+ Prod0_10[3] Prod0_10[2] Prod0_10[1] Prod0_10[0]
+ Prod0_11[3] Prod0_11[2] Prod0_11[1] Prod0_11[0]
+ Prod0_12[3] Prod0_12[2] Prod0_12[1] Prod0_12[0]
+ Prod0_13[3] Prod0_13[2] Prod0_13[1] Prod0_13[0]
+ Prod0_14[3] Prod0_14[2] Prod0_14[1] Prod0_14[0]
+ Prod0_15[3] Prod0_15[2] Prod0_15[1] Prod0_15[0]
+ Prod0_16[3] Prod0_16[2] Prod0_16[1] Prod0_16[0]
+ Prod0_17[3] Prod0_17[2] Prod0_17[1] Prod0_17[0]
+ Prod0_18[3] Prod0_18[2] Prod0_18[1] Prod0_18[0]
+ Prod0_19[3] Prod0_19[2] Prod0_19[1] Prod0_19[0]
+ Prod0_20[3] Prod0_20[2] Prod0_20[1] Prod0_20[0]
+ Prod0_21[3] Prod0_21[2] Prod0_21[1] Prod0_21[0]
+ Prod0_22[3] Prod0_22[2] Prod0_22[1] Prod0_22[0]
+ Prod0_23[3] Prod0_23[2] Prod0_23[1] Prod0_23[0]
+ Prod0_24[3] Prod0_24[2] Prod0_24[1] Prod0_24[0]
+ Prod0_25[3] Prod0_25[2] Prod0_25[1] Prod0_25[0]
+ Prod0_26[3] Prod0_26[2] Prod0_26[1] Prod0_26[0]
+ Prod0_27[3] Prod0_27[2] Prod0_27[1] Prod0_27[0]
+ Prod0_28[3] Prod0_28[2] Prod0_28[1] Prod0_28[0]
+ Prod0_29[3] Prod0_29[2] Prod0_29[1] Prod0_29[0]
+ Prod0_30[3] Prod0_30[2] Prod0_30[1] Prod0_30[0]
+ Prod0_31[3] Prod0_31[2] Prod0_31[1] Prod0_31[0]
+ CIM_Wcol

X_Wcol1 in0_b in1_b in2_b in3_b in4_b in5_b in6_b in7_b in8_b in9_b
+ in10_b in11_b in12_b in13_b in14_b in15_b in16_b in17_b in18_b in19_b
+ in20_b in21_b in22_b in23_b in24_b in25_b in26_b in27_b in28_b in29_b
+ in30_b in31_b
+ Prod1_0[3] Prod1_0[2] Prod1_0[1] Prod1_0[0]
+ Prod1_1[3] Prod1_1[2] Prod1_1[1] Prod1_1[0]
+ Prod1_2[3] Prod1_2[2] Prod1_2[1] Prod1_2[0]
+ Prod1_3[3] Prod1_3[2] Prod1_3[1] Prod1_3[0]
+ Prod1_4[3] Prod1_4[2] Prod1_4[1] Prod1_4[0]
+ Prod1_5[3] Prod1_5[2] Prod1_5[1] Prod1_5[0]
+ Prod1_6[3] Prod1_6[2] Prod1_6[1] Prod1_6[0]
+ Prod1_7[3] Prod1_7[2] Prod1_7[1] Prod1_7[0]
+ Prod1_8[3] Prod1_8[2] Prod1_8[1] Prod1_8[0]
+ Prod1_9[3] Prod1_9[2] Prod1_9[1] Prod1_9[0]
+ Prod1_10[3] Prod1_10[2] Prod1_10[1] Prod1_10[0]
+ Prod1_11[3] Prod1_11[2] Prod1_11[1] Prod1_11[0]
+ Prod1_12[3] Prod1_12[2] Prod1_12[1] Prod1_12[0]
+ Prod1_13[3] Prod1_13[2] Prod1_13[1] Prod1_13[0]
+ Prod1_14[3] Prod1_14[2] Prod1_14[1] Prod1_14[0]
+ Prod1_15[3] Prod1_15[2] Prod1_15[1] Prod1_15[0]
+ Prod1_16[3] Prod1_16[2] Prod1_16[1] Prod1_16[0]
+ Prod1_17[3] Prod1_17[2] Prod1_17[1] Prod1_17[0]
+ Prod1_18[3] Prod1_18[2] Prod1_18[1] Prod1_18[0]
+ Prod1_19[3] Prod1_19[2] Prod1_19[1] Prod1_19[0]
+ Prod1_20[3] Prod1_20[2] Prod1_20[1] Prod1_20[0]
+ Prod1_21[3] Prod1_21[2] Prod1_21[1] Prod1_21[0]
+ Prod1_22[3] Prod1_22[2] Prod1_22[1] Prod1_22[0]
+ Prod1_23[3] Prod1_23[2] Prod1_23[1] Prod1_23[0]
+ Prod1_24[3] Prod1_24[2] Prod1_24[1] Prod1_24[0]
+ Prod1_25[3] Prod1_25[2] Prod1_25[1] Prod1_25[0]
+ Prod1_26[3] Prod1_26[2] Prod1_26[1] Prod1_26[0]
+ Prod1_27[3] Prod1_27[2] Prod1_27[1] Prod1_27[0]
+ Prod1_28[3] Prod1_28[2] Prod1_28[1] Prod1_28[0]
+ Prod1_29[3] Prod1_29[2] Prod1_29[1] Prod1_29[0]
+ Prod1_30[3] Prod1_30[2] Prod1_30[1] Prod1_30[0]
+ Prod1_31[3] Prod1_31[2] Prod1_31[1] Prod1_31[0]
+ CIM_Wcol

X_Wcol2 in0_b in1_b in2_b in3_b in4_b in5_b in6_b in7_b in8_b in9_b
+ in10_b in11_b in12_b in13_b in14_b in15_b in16_b in17_b in18_b in19_b
+ in20_b in21_b in22_b in23_b in24_b in25_b in26_b in27_b in28_b in29_b
+ in30_b in31_b
+ Prod2_0[3] Prod2_0[2] Prod2_0[1] Prod2_0[0]
+ Prod2_1[3] Prod2_1[2] Prod2_1[1] Prod2_1[0]
+ Prod2_2[3] Prod2_2[2] Prod2_2[1] Prod2_2[0]
+ Prod2_3[3] Prod2_3[2] Prod2_3[1] Prod2_3[0]
+ Prod2_4[3] Prod2_4[2] Prod2_4[1] Prod2_4[0]
+ Prod2_5[3] Prod2_5[2] Prod2_5[1] Prod2_5[0]
+ Prod2_6[3] Prod2_6[2] Prod2_6[1] Prod2_6[0]
+ Prod2_7[3] Prod2_7[2] Prod2_7[1] Prod2_7[0]
+ Prod2_8[3] Prod2_8[2] Prod2_8[1] Prod2_8[0]
+ Prod2_9[3] Prod2_9[2] Prod2_9[1] Prod2_9[0]
+ Prod2_10[3] Prod2_10[2] Prod2_10[1] Prod2_10[0]
+ Prod2_11[3] Prod2_11[2] Prod2_11[1] Prod2_11[0]
+ Prod2_12[3] Prod2_12[2] Prod2_12[1] Prod2_12[0]
+ Prod2_13[3] Prod2_13[2] Prod2_13[1] Prod2_13[0]
+ Prod2_14[3] Prod2_14[2] Prod2_14[1] Prod2_14[0]
+ Prod2_15[3] Prod2_15[2] Prod2_15[1] Prod2_15[0]
+ Prod2_16[3] Prod2_16[2] Prod2_16[1] Prod2_16[0]
+ Prod2_17[3] Prod2_17[2] Prod2_17[1] Prod2_17[0]
+ Prod2_18[3] Prod2_18[2] Prod2_18[1] Prod2_18[0]
+ Prod2_19[3] Prod2_19[2] Prod2_19[1] Prod2_19[0]
+ Prod2_20[3] Prod2_20[2] Prod2_20[1] Prod2_20[0]
+ Prod2_21[3] Prod2_21[2] Prod2_21[1] Prod2_21[0]
+ Prod2_22[3] Prod2_22[2] Prod2_22[1] Prod2_22[0]
+ Prod2_23[3] Prod2_23[2] Prod2_23[1] Prod2_23[0]
+ Prod2_24[3] Prod2_24[2] Prod2_24[1] Prod2_24[0]
+ Prod2_25[3] Prod2_25[2] Prod2_25[1] Prod2_25[0]
+ Prod2_26[3] Prod2_26[2] Prod2_26[1] Prod2_26[0]
+ Prod2_27[3] Prod2_27[2] Prod2_27[1] Prod2_27[0]
+ Prod2_28[3] Prod2_28[2] Prod2_28[1] Prod2_28[0]
+ Prod2_29[3] Prod2_29[2] Prod2_29[1] Prod2_29[0]
+ Prod2_30[3] Prod2_30[2] Prod2_30[1] Prod2_30[0]
+ Prod2_31[3] Prod2_31[2] Prod2_31[1] Prod2_31[0]
+ CIM_Wcol

X_Wcol3 in0_b in1_b in2_b in3_b in4_b in5_b in6_b in7_b in8_b in9_b
+ in10_b in11_b in12_b in13_b in14_b in15_b in16_b in17_b in18_b in19_b
+ in20_b in21_b in22_b in23_b in24_b in25_b in26_b in27_b in28_b in29_b
+ in30_b in31_b
+ Prod3_0[3] Prod3_0[2] Prod3_0[1] Prod3_0[0]
+ Prod3_1[3] Prod3_1[2] Prod3_1[1] Prod3_1[0]
+ Prod3_2[3] Prod3_2[2] Prod3_2[1] Prod3_2[0]
+ Prod3_3[3] Prod3_3[2] Prod3_3[1] Prod3_3[0]
+ Prod3_4[3] Prod3_4[2] Prod3_4[1] Prod3_4[0]
+ Prod3_5[3] Prod3_5[2] Prod3_5[1] Prod3_5[0]
+ Prod3_6[3] Prod3_6[2] Prod3_6[1] Prod3_6[0]
+ Prod3_7[3] Prod3_7[2] Prod3_7[1] Prod3_7[0]
+ Prod3_8[3] Prod3_8[2] Prod3_8[1] Prod3_8[0]
+ Prod3_9[3] Prod3_9[2] Prod3_9[1] Prod3_9[0]
+ Prod3_10[3] Prod3_10[2] Prod3_10[1] Prod3_10[0]
+ Prod3_11[3] Prod3_11[2] Prod3_11[1] Prod3_11[0]
+ Prod3_12[3] Prod3_12[2] Prod3_12[1] Prod3_12[0]
+ Prod3_13[3] Prod3_13[2] Prod3_13[1] Prod3_13[0]
+ Prod3_14[3] Prod3_14[2] Prod3_14[1] Prod3_14[0]
+ Prod3_15[3] Prod3_15[2] Prod3_15[1] Prod3_15[0]
+ Prod3_16[3] Prod3_16[2] Prod3_16[1] Prod3_16[0]
+ Prod3_17[3] Prod3_17[2] Prod3_17[1] Prod3_17[0]
+ Prod3_18[3] Prod3_18[2] Prod3_18[1] Prod3_18[0]
+ Prod3_19[3] Prod3_19[2] Prod3_19[1] Prod3_19[0]
+ Prod3_20[3] Prod3_20[2] Prod3_20[1] Prod3_20[0]
+ Prod3_21[3] Prod3_21[2] Prod3_21[1] Prod3_21[0]
+ Prod3_22[3] Prod3_22[2] Prod3_22[1] Prod3_22[0]
+ Prod3_23[3] Prod3_23[2] Prod3_23[1] Prod3_23[0]
+ Prod3_24[3] Prod3_24[2] Prod3_24[1] Prod3_24[0]
+ Prod3_25[3] Prod3_25[2] Prod3_25[1] Prod3_25[0]
+ Prod3_26[3] Prod3_26[2] Prod3_26[1] Prod3_26[0]
+ Prod3_27[3] Prod3_27[2] Prod3_27[1] Prod3_27[0]
+ Prod3_28[3] Prod3_28[2] Prod3_28[1] Prod3_28[0]
+ Prod3_29[3] Prod3_29[2] Prod3_29[1] Prod3_29[0]
+ Prod3_30[3] Prod3_30[2] Prod3_30[1] Prod3_30[0]
+ Prod3_31[3] Prod3_31[2] Prod3_31[1] Prod3_31[0]
+ CIM_Wcol
.ends

.subckt CIM_Wcol
+ in0_b in1_b in2_b in3_b in4_b in5_b in6_b in7_b in8_b in9_b
+ in10_b in11_b in12_b in13_b in14_b in15_b in16_b in17_b in18_b in19_b
+ in20_b in21_b in22_b in23_b in24_b in25_b in26_b in27_b in28_b in29_b
+ in30_b in31_b
+ Prod0[3] Prod0[2] Prod0[1] Prod0[0]
+ Prod1[3] Prod1[2] Prod1[1] Prod1[0]
+ Prod2[3] Prod2[2] Prod2[1] Prod2[0]
+ Prod3[3] Prod3[2] Prod3[1] Prod3[0]
+ Prod4[3] Prod4[2] Prod4[1] Prod4[0]
+ Prod5[3] Prod5[2] Prod5[1] Prod5[0]
+ Prod6[3] Prod6[2] Prod6[1] Prod6[0]
+ Prod7[3] Prod7[2] Prod7[1] Prod7[0]
+ Prod8[3] Prod8[2] Prod8[1] Prod8[0]
+ Prod9[3] Prod9[2] Prod9[1] Prod9[0]
+ Prod10[3] Prod10[2] Prod10[1] Prod10[0]
+ Prod11[3] Prod11[2] Prod11[1] Prod11[0]
+ Prod12[3] Prod12[2] Prod12[1] Prod12[0]
+ Prod13[3] Prod13[2] Prod13[1] Prod13[0]
+ Prod14[3] Prod14[2] Prod14[1] Prod14[0]
+ Prod15[3] Prod15[2] Prod15[1] Prod15[0]
+ Prod16[3] Prod16[2] Prod16[1] Prod16[0]
+ Prod17[3] Prod17[2] Prod17[1] Prod17[0]
+ Prod18[3] Prod18[2] Prod18[1] Prod18[0]
+ Prod19[3] Prod19[2] Prod19[1] Prod19[0]
+ Prod20[3] Prod20[2] Prod20[1] Prod20[0]
+ Prod21[3] Prod21[2] Prod21[1] Prod21[0]
+ Prod22[3] Prod22[2] Prod22[1] Prod22[0]
+ Prod23[3] Prod23[2] Prod23[1] Prod23[0]
+ Prod24[3] Prod24[2] Prod24[1] Prod24[0]
+ Prod25[3] Prod25[2] Prod25[1] Prod25[0]
+ Prod26[3] Prod26[2] Prod26[1] Prod26[0]
+ Prod27[3] Prod27[2] Prod27[1] Prod27[0]
+ Prod28[3] Prod28[2] Prod28[1] Prod28[0]
+ Prod29[3] Prod29[2] Prod29[1] Prod29[0]
+ Prod30[3] Prod30[2] Prod30[1] Prod30[0]
+ Prod31[3] Prod31[2] Prod31[1] Prod31[0]


X_W0 in0_b Prod0[3] Prod0[2] Prod0[1] Prod0[0] CIM_W
X_W1 in1_b Prod1[3] Prod1[2] Prod1[1] Prod1[0] CIM_W
X_W2 in2_b Prod2[3] Prod2[2] Prod2[1] Prod2[0] CIM_W
X_W3 in3_b Prod3[3] Prod3[2] Prod3[1] Prod3[0] CIM_W
X_W4 in4_b Prod4[3] Prod4[2] Prod4[1] Prod4[0] CIM_W
X_W5 in5_b Prod5[3] Prod5[2] Prod5[1] Prod5[0] CIM_W
X_W6 in6_b Prod6[3] Prod6[2] Prod6[1] Prod6[0] CIM_W
X_W7 in7_b Prod7[3] Prod7[2] Prod7[1] Prod7[0] CIM_W
X_W8 in8_b Prod8[3] Prod8[2] Prod8[1] Prod8[0] CIM_W
X_W9 in9_b Prod9[3] Prod9[2] Prod9[1] Prod9[0] CIM_W

X_W10 in10_b Prod10[3] Prod10[2] Prod10[1] Prod10[0] CIM_W
X_W11 in11_b Prod11[3] Prod11[2] Prod11[1] Prod11[0] CIM_W
X_W12 in12_b Prod12[3] Prod12[2] Prod12[1] Prod12[0] CIM_W
X_W13 in13_b Prod13[3] Prod13[2] Prod13[1] Prod13[0] CIM_W
X_W14 in14_b Prod14[3] Prod14[2] Prod14[1] Prod14[0] CIM_W
X_W15 in15_b Prod15[3] Prod15[2] Prod15[1] Prod15[0] CIM_W
X_W16 in16_b Prod16[3] Prod16[2] Prod16[1] Prod16[0] CIM_W
X_W17 in17_b Prod17[3] Prod17[2] Prod17[1] Prod17[0] CIM_W
X_W18 in18_b Prod18[3] Prod18[2] Prod18[1] Prod18[0] CIM_W
X_W19 in19_b Prod19[3] Prod19[2] Prod19[1] Prod19[0] CIM_W

X_W20 in20_b Prod20[3] Prod20[2] Prod20[1] Prod20[0] CIM_W
X_W21 in21_b Prod21[3] Prod21[2] Prod21[1] Prod21[0] CIM_W
X_W22 in22_b Prod22[3] Prod22[2] Prod22[1] Prod22[0] CIM_W
X_W23 in23_b Prod23[3] Prod23[2] Prod23[1] Prod23[0] CIM_W
X_W24 in24_b Prod24[3] Prod24[2] Prod24[1] Prod24[0] CIM_W
X_W25 in25_b Prod25[3] Prod25[2] Prod25[1] Prod25[0] CIM_W
X_W26 in26_b Prod26[3] Prod26[2] Prod26[1] Prod26[0] CIM_W
X_W27 in27_b Prod27[3] Prod27[2] Prod27[1] Prod27[0] CIM_W
X_W28 in28_b Prod28[3] Prod28[2] Prod28[1] Prod28[0] CIM_W
X_W29 in29_b Prod29[3] Prod29[2] Prod29[1] Prod29[0] CIM_W

X_W30 in30_b Prod30[3] Prod30[2] Prod30[1] Prod30[0] CIM_W
X_W31 in31_b Prod31[3] Prod31[2] Prod31[1] Prod31[0] CIM_W
.ends

.subckt CIM_W I P[3] P[2] P[1] P[0]
X_bit0 I P[0] WL[0] BL[0] BLB[0] W[0] qb[0] CIM_cell
X_bit1 I P[1] WL[0] BL[1] BLB[1] W[1] qb[1] CIM_cell
X_bit2 I P[2] WL[0] BL[2] BLB[2] W[2] qb[2] CIM_cell
X_bit3 I P[3] WL[0] BL[3] BLB[3] W[3] qb[3] CIM_cell
.IC V(BL[0]) = 0V
.IC V(BL[1]) = 0V
.IC V(BL[2]) = 0V
.IC V(BL[3]) = 0V
.IC V(BLB[0]) = 0V
.IC V(BLB[1]) = 0V
.IC V(BLB[2]) = 0V
.IC V(BLB[3]) = 0V 
.IC V(WL[0]) = 0V
.ends

