.SUBCKT Accumulators VPRW VGND  rst_n clk
+ P[8] P[7] P[6] P[5] P[4] P[3] P[2] P[1] P[0]
+ out_valid O[12] O[11] O[10] O[9] O[8] O[7] O[6] O[5] O[4] O[3] O[2] O[1] O[0]
XU84 ctr[0] n151 ctr[1] ctr[4] ctr[2] VPRW VGND  N57 NOR5xp2_ASAP7_75t_R
XU95 N7 n72 VPRW VGND  n76 AND2x2_ASAP7_75t_R
XU96 ctr[1] n151 flag VPRW VGND  n75 AND3x1_ASAP7_75t_R
Xadd_63 VPRW VGND  n1 n1 n1 n1 P[8] P[7] P[6] P[5] P[4] P[3] P[2] P[1] P[0]
+ O[11] O[10] O[9] O[8] O[7] O[6] O[5] O[4] O[3] O[2] O[1] O[0]
+ n1 n1 N43 N42 N41 N40 N39 N38 N37 N36 N35 N34 N33 N32 N31 CO_f1
+ Accumulators_DW01_add_0
*.SUBCKT HAxp5_ASAP7_75t_R A B CON SN VDD VSS
Xadd_39_U1_1_1 ctr[1] ctr[0] n128 n127 VPRW VGND HAxp5_ASAP7_75t_R
Xadd_39_U1_1_2 ctr[2] n133 n130 n129 VPRW VGND HAxp5_ASAP7_75t_R
Xadd_39_U1_1_3 ctr[3] n134 n132 n131 VPRW VGND HAxp5_ASAP7_75t_R
Xflag_reg clk n83 flag n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg clk n82 out_valid n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
Xctr_reg_2_ clk n81 ctr[2] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
Xctr_reg_1_ clk n80 ctr[1] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
Xctr_reg_0_ clk n79 ctr[0] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
Xctr_reg_3_ clk n77 ctr[3] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
Xctr_reg_4_ clk n78 ctr[4] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_0_ clk n150 O[0] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_1_ clk n149 O[1] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_2_ clk n148 O[2] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_3_ clk n147 O[3] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_4_ clk n146 O[4] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_5_ clk n145 O[5] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_6_ clk n144 O[6] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_7_ clk n143 O[7] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_8_ clk n142 O[8] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_11_ clk n139 O[11] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_12_ clk n138 O[12] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_10_ clk n140 O[10] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XO_reg_9_ clk n141 O[9] n126 n1 VPRW VGND ASYNC_DFFHx1_ASAP7_75t_R
XU97 n1 VPRW VGND  TIELOx1_ASAP7_75t_R
XU98 n125 N43 VPRW VGND  n138 NAND2xp5_ASAP7_75t_R
XU99 N14 n76 VPRW VGND  n77 NAND2xp5_ASAP7_75t_R
XU100 N15 n76 VPRW VGND  n78 NAND2xp5_ASAP7_75t_R
XU101 N11 n76 VPRW VGND  n79 NAND2xp5_ASAP7_75t_R
XU102 N12 n76 VPRW VGND  n80 NAND2xp5_ASAP7_75t_R
XU103 N13 n76 VPRW VGND  n81 NAND2xp5_ASAP7_75t_R
XU104 ctr[4] ctr[2] ctr[0] n73 VPRW VGND  n82 OR4x2_ASAP7_75t_R
XU105 flag N57 VPRW VGND  n83 NOR2xp33_ASAP7_75t_R
XU106 n122 VPRW VGND  n125 INVx1_ASAP7_75t_R
XU107 n87 n72 VPRW VGND  n122 NAND2xp5_ASAP7_75t_R
XU108 ctr[3] ctr[0] n86 n85 VPRW VGND  n87 NAND4xp25_ASAP7_75t_R
XU109 ctr[1] ctr[2] VPRW VGND  n85 NOR2xp33_ASAP7_75t_R
XU110 ctr[2] ctr[4] VPRW VGND  n84 NOR2xp33_ASAP7_75t_R
XU111 n74 n75 VPRW VGND  n73 NOR2xp33_ASAP7_75t_R
XU112 ctr[1] n151 VPRW VGND  n74 NOR2xp33_ASAP7_75t_R
XU113 n75 ctr[0] n84 VPRW VGND  n72 NAND3xp33_ASAP7_75t_R
XU114 rst_n VPRW VGND  n126 INVx1_ASAP7_75t_R
XU115 ctr[4] VPRW VGND  n86 INVx1_ASAP7_75t_R
XU116 N42 n125 VPRW VGND  n139 NAND2xp5_ASAP7_75t_R
XU117 N41 n125 VPRW VGND  n140 NAND2xp5_ASAP7_75t_R
XU118 N40 n125 VPRW VGND  n141 NAND2xp5_ASAP7_75t_R
XU119 N39 VPRW VGND  n88 INVx1_ASAP7_75t_R
XU120 n125 n88 VPRW VGND  n91 NAND2xp5_ASAP7_75t_R
XU121 P[8] VPRW VGND  n89 INVx1_ASAP7_75t_R
XU122 n122 n89 VPRW VGND  n90 NAND2xp5_ASAP7_75t_R
XU123 n91 n90 VPRW VGND  n142 NAND2xp5_ASAP7_75t_R
XU124 N38 VPRW VGND  n92 INVx1_ASAP7_75t_R
XU125 n125 n92 VPRW VGND  n95 NAND2xp5_ASAP7_75t_R
XU126 P[7] VPRW VGND  n93 INVx1_ASAP7_75t_R
XU127 n122 n93 VPRW VGND  n94 NAND2xp5_ASAP7_75t_R
XU128 n95 n94 VPRW VGND  n143 NAND2xp5_ASAP7_75t_R
XU129 N37 VPRW VGND  n96 INVx1_ASAP7_75t_R
XU130 n125 n96 VPRW VGND  n99 NAND2xp5_ASAP7_75t_R
XU131 P[6] VPRW VGND  n97 INVx1_ASAP7_75t_R
XU132 n122 n97 VPRW VGND  n98 NAND2xp5_ASAP7_75t_R
XU133 n99 n98 VPRW VGND  n144 NAND2xp5_ASAP7_75t_R
XU134 N36 VPRW VGND  n100 INVx1_ASAP7_75t_R
XU135 n125 n100 VPRW VGND  n103 NAND2xp5_ASAP7_75t_R
XU136 P[5] VPRW VGND  n101 INVx1_ASAP7_75t_R
XU137 n122 n101 VPRW VGND  n102 NAND2xp5_ASAP7_75t_R
XU138 n103 n102 VPRW VGND  n145 NAND2xp5_ASAP7_75t_R
XU139 N35 VPRW VGND  n104 INVx1_ASAP7_75t_R
XU140 n125 n104 VPRW VGND  n107 NAND2xp5_ASAP7_75t_R
XU141 P[4] VPRW VGND  n105 INVx1_ASAP7_75t_R
XU142 n122 n105 VPRW VGND  n106 NAND2xp5_ASAP7_75t_R
XU143 n107 n106 VPRW VGND  n146 NAND2xp5_ASAP7_75t_R
XU144 N34 VPRW VGND  n108 INVx1_ASAP7_75t_R
XU145 n125 n108 VPRW VGND  n111 NAND2xp5_ASAP7_75t_R
XU146 P[3] VPRW VGND  n109 INVx1_ASAP7_75t_R
XU147 n122 n109 VPRW VGND  n110 NAND2xp5_ASAP7_75t_R
XU148 n111 n110 VPRW VGND  n147 NAND2xp5_ASAP7_75t_R
XU149 N33 VPRW VGND  n112 INVx1_ASAP7_75t_R
XU150 n125 n112 VPRW VGND  n115 NAND2xp5_ASAP7_75t_R
XU151 P[2] VPRW VGND  n113 INVx1_ASAP7_75t_R
XU152 n122 n113 VPRW VGND  n114 NAND2xp5_ASAP7_75t_R
XU153 n115 n114 VPRW VGND  n148 NAND2xp5_ASAP7_75t_R
XU154 N32 VPRW VGND  n116 INVx1_ASAP7_75t_R
XU155 n125 n116 VPRW VGND  n119 NAND2xp5_ASAP7_75t_R
XU156 P[1] VPRW VGND  n117 INVx1_ASAP7_75t_R
XU157 n122 n117 VPRW VGND  n118 NAND2xp5_ASAP7_75t_R
XU158 n119 n118 VPRW VGND  n149 NAND2xp5_ASAP7_75t_R
XU159 N31 VPRW VGND  n120 INVx1_ASAP7_75t_R
XU160 n125 n120 VPRW VGND  n124 NAND2xp5_ASAP7_75t_R
XU161 P[0] VPRW VGND  n121 INVx1_ASAP7_75t_R
XU162 n122 n121 VPRW VGND  n123 NAND2xp5_ASAP7_75t_R
XU163 n124 n123 VPRW VGND  n150 NAND2xp5_ASAP7_75t_R
XU164 ctr[0] VPRW VGND  N11 INVx1_ASAP7_75t_R
XU165 n127 VPRW VGND  N12 INVx1_ASAP7_75t_R
XU166 n129 VPRW VGND  N13 INVx1_ASAP7_75t_R
XU167 n131 VPRW VGND  N14 INVx1_ASAP7_75t_R
XU168 n132 ctr[4] VPRW VGND  N15 XNOR2xp5_ASAP7_75t_R
XU169 n128 VPRW VGND  n133 INVx1_ASAP7_75t_R
XU170 n130 VPRW VGND  n134 INVx1_ASAP7_75t_R
XU171 ctr[0] ctr[1] VPRW VGND  n135 NOR2xp33_ASAP7_75t_R
XU172 n135 n151 VPRW VGND  n137 NOR2xp33_ASAP7_75t_R
XU173 ctr[3] ctr[2] VPRW VGND  n136 AND2x2_ASAP7_75t_R
XU174 n137 ctr[4] n136 VPRW VGND  N7 NOR3xp33_ASAP7_75t_R
XU175 ctr[3] VPRW VGND  n151 INVx1_ASAP7_75t_R
.ENDS




