.SUBCKT Adder_Tree_DW01_add_5 VPRW VGND  A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_5 A[5] B[5] n3 n7 n8  VPRW VGND  FAx1_ASAP7_75t_R
XU1_4 A[4] B[4] n4 n9 n10  VPRW VGND  FAx1_ASAP7_75t_R
XU1_3 A[3] B[3] n5 n11 n12  VPRW VGND  FAx1_ASAP7_75t_R
XU1_2 A[2] B[2] n6 n13 n14  VPRW VGND  FAx1_ASAP7_75t_R
XU1_1 A[1] B[1] n1 n15 n16  VPRW VGND  FAx1_ASAP7_75t_R
XU1 A[0] B[0] VPRW VGND  n1 AND2x2_ASAP7_75t_R
XU2 B[0] A[0] VPRW VGND  SUM[0] XOR2xp5_ASAP7_75t_R
XU3 n9 VPRW VGND  n3 INVx1_ASAP7_75t_R
XU4 n11 VPRW VGND  n4 INVx1_ASAP7_75t_R
XU5 n13 VPRW VGND  n5 INVx1_ASAP7_75t_R
XU6 n15 VPRW VGND  n6 INVx1_ASAP7_75t_R
XU7 n7 VPRW VGND  SUM[6] INVx1_ASAP7_75t_R
XU8 n8 VPRW VGND  SUM[5] INVx1_ASAP7_75t_R
XU9 n10 VPRW VGND  SUM[4] INVx1_ASAP7_75t_R
XU10 n12 VPRW VGND  SUM[3] INVx1_ASAP7_75t_R
XU11 n14 VPRW VGND  SUM[2] INVx1_ASAP7_75t_R
XU12 n16 VPRW VGND  SUM[1] INVx1_ASAP7_75t_R
.ENDS


