.SUBCKT Accumulators_DW01_add_0 VPRW VGND  A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_8 A[8] B[8] n15 n22 n23  VPRW VGND  FAx1_ASAP7_75t_R
XU1_7 A[7] B[7] n16 n24 n25  VPRW VGND  FAx1_ASAP7_75t_R
XU1_6 A[6] B[6] n17 n26 n27  VPRW VGND  FAx1_ASAP7_75t_R
XU1_5 A[5] B[5] n18 n28 n29  VPRW VGND  FAx1_ASAP7_75t_R
XU1_4 A[4] B[4] n19 n30 n31  VPRW VGND  FAx1_ASAP7_75t_R
XU1_3 A[3] B[3] n20 n32 n33  VPRW VGND  FAx1_ASAP7_75t_R
XU1_2 A[2] B[2] n7 n34 n35  VPRW VGND  FAx1_ASAP7_75t_R
XU1 n22 n2 VPRW VGND  n9 NOR2xp33_ASAP7_75t_R
XU2 B[9] B[10] VPRW VGND  n2 NAND2xp5_ASAP7_75t_R
XU3 n8 B[10] VPRW VGND  SUM[10] XOR2xp5_ASAP7_75t_R
XU4 B[11] n9 VPRW VGND  n21 NAND2xp5_ASAP7_75t_R
XU5 B[11] VPRW VGND  n4 INVx1_ASAP7_75t_R
XU6 n14 B[9] VPRW VGND  SUM[9] XOR2xp5_ASAP7_75t_R
XU7 n9 n4 VPRW VGND  SUM[11] XNOR2xp5_ASAP7_75t_R
XU8 A[1] VPRW VGND  n5 INVx8_ASAP7_75t_R
XU9 n5 n6 VPRW VGND  n7 NOR2x1p5_ASAP7_75t_R
XU10 B[1] VPRW VGND  n6 INVx13_ASAP7_75t_R
XU11 B[9] n14 VPRW VGND  n8 AND2x2_ASAP7_75t_R
XU12 n21 B[12] VPRW VGND  SUM[12] XNOR2xp5_ASAP7_75t_R
XU13 B[1] A[1] VPRW VGND  SUM[1] XOR2xp5_ASAP7_75t_R
XU14 A[0] VPRW VGND  SUM[0] HB1xp67_ASAP7_75t_R
XU15 n22 VPRW VGND  n14 INVx1_ASAP7_75t_R
XU16 n24 VPRW VGND  n15 INVx1_ASAP7_75t_R
XU17 n26 VPRW VGND  n16 INVx1_ASAP7_75t_R
XU18 n28 VPRW VGND  n17 INVx1_ASAP7_75t_R
XU19 n30 VPRW VGND  n18 INVx1_ASAP7_75t_R
XU20 n32 VPRW VGND  n19 INVx1_ASAP7_75t_R
XU21 n34 VPRW VGND  n20 INVx1_ASAP7_75t_R
XU22 n23 VPRW VGND  SUM[8] INVx1_ASAP7_75t_R
XU23 n25 VPRW VGND  SUM[7] INVx1_ASAP7_75t_R
XU24 n27 VPRW VGND  SUM[6] INVx1_ASAP7_75t_R
XU25 n29 VPRW VGND  SUM[5] INVx1_ASAP7_75t_R
XU26 n31 VPRW VGND  SUM[4] INVx1_ASAP7_75t_R
XU27 n33 VPRW VGND  SUM[3] INVx1_ASAP7_75t_R
XU28 n35 VPRW VGND  SUM[2] INVx1_ASAP7_75t_R
.ENDS

