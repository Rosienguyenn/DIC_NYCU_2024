
.subckt buffer_arr 
+ a[0] y[0] a[1] y[1] a[2] y[2] a[3] y[3] a[4] y[4]
+ a[5] y[5] a[6] y[6] a[7] y[7] a[8] y[8] a[9] y[9]
+ a[10] y[10] a[11] y[11] a[12] y[12] a[13] y[13] a[14] y[14]
+ a[15] y[15] a[16] y[16] a[17] y[17] a[18] y[18] a[19] y[19]
+ a[20] y[20] a[21] y[21] a[22] y[22] a[23] y[23] a[24] y[24]
+ a[25] y[25] a[26] y[26] a[27] y[27] a[28] y[28] a[29] y[29]
+ a[30] y[30] a[31] y[31]

x_buf0 a[0] y[0] Buffer
x_buf1 a[1] y[1] Buffer
x_buf2 a[2] y[2] Buffer
x_buf3 a[3] y[3] Buffer
x_buf4 a[4] y[4] Buffer
x_buf5 a[5] y[5] Buffer
x_buf6 a[6] y[6] Buffer
x_buf7 a[7] y[7] Buffer
x_buf8 a[8] y[8] Buffer
x_buf9 a[9] y[9] Buffer

x_buf10 a[10] y[10] Buffer
x_buf11 a[11] y[11] Buffer
x_buf12 a[12] y[12] Buffer
x_buf13 a[13] y[13] Buffer
x_buf14 a[14] y[14] Buffer
x_buf15 a[15] y[15] Buffer
x_buf16 a[16] y[16] Buffer
x_buf17 a[17] y[17] Buffer
x_buf18 a[18] y[18] Buffer
x_buf19 a[19] y[19] Buffer

x_buf20 a[20] y[20] Buffer
x_buf21 a[21] y[21] Buffer
x_buf22 a[22] y[22] Buffer
x_buf23 a[23] y[23] Buffer
x_buf24 a[24] y[24] Buffer
x_buf25 a[25] y[25] Buffer
x_buf26 a[26] y[26] Buffer
x_buf27 a[27] y[27] Buffer
x_buf28 a[28] y[28] Buffer
x_buf29 a[29] y[29] Buffer

x_buf30 a[30] y[30] Buffer
x_buf31 a[31] y[31] Buffer
.ends
